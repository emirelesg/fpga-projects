`ifndef _IO_MMIO_MAP_INCLUDED
`define _IO_MMIO_MAP_INCLUDED

// Slot definition
`define S0_LED 0

`endif
