/*
 * uart_baudrate_gen
 * 
 */

module uart_baudrate_gen
    (
        input logic clk,
        input logic reset_n
    );

endmodule
