`ifndef _IO_MMIO_MAP_INCLUDED
`define _IO_MMIO_MAP_INCLUDED

// Slot definition
`define IO_S0_GPO 0
`define IO_S1_DDFS 1

`endif
