module top
    (
        input logic clk,
        input logic reset_n
    );

endmodule
