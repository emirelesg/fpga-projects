module delay
    (
        input logic i_clk,
        input logic i_reset_n
    );

endmodule
