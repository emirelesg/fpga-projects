/*
 * uart_tx
 * 
 */

module uart_tx
    (
        input logic clk,
        input logic reset_n
    );

endmodule
