module top
    (

    );

endmodule
