`timescale 1ns / 10ps

module reg_file_tb;
    localparam T=10; // 100 Mhz, 10 ns

    logic clk;
    logic reset_n;

    localparam DATA_WIDTH = 8;
    localparam ADDR_WIDTH = 3;

    logic wr_en;
    logic [ADDR_WIDTH-1:0] wr_addr, rd_addr;
    logic [DATA_WIDTH-1:0] wr_data, rd_data;

    reg_file #(.DATA_WIDTH(DATA_WIDTH), .ADDR_WIDTH(ADDR_WIDTH)) uut(
        .clk(clk),
        .reset_n(reset_n),
        .wr_en(wr_en),
        .wr_addr(wr_addr),
        .rd_addr(rd_addr),
        .wr_data(wr_data),
        .rd_data(rd_data)
    );

    // Simulate a 100 Mhz clock signal.
    always begin
        clk = 1'b0;
        #(T/2);
        clk = 1'b1;
        #(T/2);
    end

    // Reset at the start of the simulation.
    initial begin
        wr_en = 1'b0;
        wr_addr = 2'b00;
        wr_data = 8'h00;
        rd_addr = 2'b00;

        reset_n = 1'b0;
        #(T/2);
        reset_n = 1'b1;
        #(T);
    end

    initial begin
        @(posedge reset_n); // Wait for the reset.
        @(negedge clk);

        // Write to all addresses a byte.
        wr_en = 1'b1;
        for (logic [DATA_WIDTH-1:0] i=0; i < 2**ADDR_WIDTH; i++) begin
            wr_addr = i;
            wr_data = 8'hff - i;
            @(negedge clk);
        end
        wr_en = 1'b0;
        wr_addr = 2'b00;
        wr_data = 8'h00;

        // Read all addresses.
        for (logic [DATA_WIDTH-1:0] i=0; i < 2**ADDR_WIDTH; i++) begin
            rd_addr = i;
            @(negedge clk);
        end

        $stop;
    end
endmodule
