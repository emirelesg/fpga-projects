module adsr
    (
        input logic clk,
        input logic reset_n
    );

endmodule
