module i2s
    (
        input logic clk_i2s,
        input logic reset_n
    );

endmodule
